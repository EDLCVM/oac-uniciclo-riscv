library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.riscv_pkg.all;

entity ULAControle is
	port (
		ALUOp : out ULA_OP
	);
end ULAControle;

architecture comportamento of ULAControle is
begin
end comportamento;