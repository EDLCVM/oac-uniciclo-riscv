library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.riscv_pkg.all;

entity Processador is
end Processador;

architecture comportamento of Processador is
begin
end comportamento;