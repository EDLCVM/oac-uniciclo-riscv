entity Adder is
end Adder;

architecture comportamento of Adder is
begin
end comportamento;